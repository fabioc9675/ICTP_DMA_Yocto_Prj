----------------------------------------------------------------------------------
-- Generador de medio círculo (semicircular wave)
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity semicircle_wave_gen is
    Port ( 
            clk        : in  STD_LOGIC;
            rst        : in  STD_LOGIC;
            semi_out   : out STD_LOGIC_VECTOR (15 downto 0)
         );
end semicircle_wave_gen;

architecture Behavioral of semicircle_wave_gen is

    type semicircle_table is array(0 to 255) of integer range 0 to 65535;
    constant semi_table : semicircle_table := (
     0,  8192, 11562, 14133, 16287, 18173, 19867, 21416,
 22849, 24186, 25442, 26628, 27755, 28834, 29870, 30870,
 31838, 32777, 33689, 34577, 35444, 36291, 37119, 37930,
 38724, 39504, 40269, 41021, 41760, 42487, 43203, 43909,
 44604, 45289, 45965, 46632, 47291, 47942, 48585, 49220,
 49849, 50470, 51085, 51693, 52295, 52891, 53480, 54064,
 54642, 55214, 55780, 56341, 56896, 57445, 57989, 58528,
 59062, 59590, 60113, 60631, 61143, 61651, 62154, 62651,
 63143, 63631, 64113, 64590, 65062, 65529, 65529, 65062,
 64590, 64113, 63631, 63143, 62651, 62154, 61651, 61143,
 60631, 60113, 59590, 59062, 58528, 57989, 57445, 56896,
 56341, 55780, 55214, 54642, 54064, 53480, 52891, 52295,
 51693, 51085, 50470, 49849, 49220, 48585, 47942, 47291,
 46632, 45965, 45289, 44604, 43909, 43203, 42487, 41760,
 41021, 40269, 39504, 38724, 37930, 37119, 36291, 35444,
 34577, 33689, 32777, 31838, 30870, 29870, 28834, 27755,
 26628, 25442, 24186, 22849, 21416, 19867, 18173, 16287,
 14133, 11562,  8192,     0,     0,  8192, 11562, 14133,
 16287, 18173, 19867, 21416, 22849, 24186, 25442, 26628,
 27755, 28834, 29870, 30870, 31838, 32777, 33689, 34577,
 35444, 36291, 37119, 37930, 38724, 39504, 40269, 41021,
 41760, 42487, 43203, 43909, 44604, 45289, 45965, 46632,
 47291, 47942, 48585, 49220, 49849, 50470, 51085, 51693,
 52295, 52891, 53480, 54064, 54642, 55214, 55780, 56341,
 56896, 57445, 57989, 58528, 59062, 59590, 60113, 60631,
 61143, 61651, 62154, 62651, 63143, 63631, 64113, 64590,
 65062, 65529, 65529, 65062, 64590, 64113, 63631, 63143,
 62651, 62154, 61651, 61143, 60631, 60113, 59590, 59062,
 58528, 57989, 57445, 56896, 56341, 55780, 55214, 54642,
 54064, 53480, 52891, 52295, 51693, 51085, 50470, 49849,
 49220, 48585, 47942, 47291, 46632, 45965, 45289, 44604,
 43909, 43203, 42487, 41760, 41021, 40269, 39504, 38724,
 37930, 37119, 36291, 35444, 34577, 33689, 32777, 31838,
 30870, 29870, 28834, 27755, 26628, 25442, 24186, 22849,
 21416, 19867, 18173, 16287, 14133, 11562,  8192,     0
);

    signal idx  : integer range 0 to 255 := 0;
    signal val  : integer range 0 to 65535 := 0;

begin
    process(clk, rst)
    begin
        if rst = '1' then
            idx <= 0;
            val <= semi_table(0);
        elsif rising_edge(clk) then
            val <= semi_table(idx);
            semi_out <= conv_std_logic_vector(val, 16);

            if idx = 255 then
                idx <= 0;
            else
                idx <= idx + 1;
            end if;
        end if;
    end process;
end Behavioral;